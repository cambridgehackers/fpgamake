
// Permission is hereby granted, free of charge, to any person
// obtaining a copy of this software and associated documentation
// files (the "Software"), to deal in the Software without
// restriction, including without limitation the rights to use, copy,
// modify, merge, publish, distribute, sublicense, and/or sell copies
// of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be
// included in all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
// EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS
// BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN
// ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN
// CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.

interface MetaHarden#(type a);
   (* always_ready, always_enabled *)
   method Action signal(a src);
   (* always_ready *)
   method a signal_dst;
endinterface
   
module mkMetaHarden#(a initVal)(MetaHarden#(a))
   provisos(Bits#(a, sa));

   Reg#(a) signal_meta <- mkReg(initVal);
   Reg#(a) signal_out  <- mkReg(initVal);
   
   rule meta_hardner;
      signal_out <= signal_meta;
   endrule
   
   method Action signal(a src);
      signal_meta <= src;
   endmethod
   
   method signal_dst = signal_out;
   
endmodule